module imm_gen(
    input [31:0] inst,
  	output reg [31:0] imm
);


    always @ (*)
        case(inst[6:0])

            7'b0000011,
          	7'b0010011:
              imm = {{20{inst[31]}}, inst[31:20]}; // lw and addi

            7'b0100011:

          		imm = {{20{inst[31]}}, inst[31:25], inst[11:7]};
          		

            7'b1100011:
      
  		 		imm = {{19{inst[31]}}, inst[7], inst[30:25], inst[11:8], 1'b0};

        endcase

endmodule

//VERIFY AND EDIT
//FINISH SIGN EXTENDING
